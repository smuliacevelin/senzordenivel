** Profile: "SCHEMATIC1-temperatura"  [ c:\users\evelin\documents\facultate\an 2 sem 2\cad\senzor_de_nivel_nou-pspicefiles\senzor_de_nivel_nou-PSpiceFiles\SCHEMATIC1\temperatura.sim ] 

** Creating circuit file "temperatura.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../leduri/red_led.lib" 
.LIB "../../../leduri/blue_led.lib" 
.LIB "../../../leduri/green_led.lib" 
.LIB "../../../leduri/yellow_led.lib" 
* From [PSPICE NETLIST] section of C:\SPB_DATA\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
